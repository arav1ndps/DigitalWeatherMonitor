library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.NUMERIC_STD.ALL;

entity alarm_tb is
end alarm_tb;

architecture arch_alarm_tb of alarm_tb is

begin


end arch_alarm_tb;
